// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_SB_ST_CHKR_SV__
`define __UVME_SB_ST_CHKR_SV__


/**
 * TODO Describe uvme_sb_st_chkr
 */
module uvme_sb_st_chkr (
      uvma_sb_if  abc_if,
      uvma_sb_if  def_if
);
   
   `pragma protect begin
   
   // TODO Add assertions to uvme_sb_st_chkr
   
   `pragma protect end
   
endmodule : uvme_sb_st_chkr


`endif // __UVME_SB_ST_CHKR_SV__
