// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_SB_MACROS_SV__
`define __UVML_SB_MACROS_SV__


`ifndef UVML_SB_MDUPLEX_MAX_CHANNELS
   `define UVML_SB_MDUPLEX_MAX_CHANNELS 8
`endif

`ifndef UVML_SB_MSIMPLEX_MAX_STREAMS
   `define UVML_SB_MSIMPLEX_MAX_STREAMS 8
`endif


`endif // __UVML_SB_MACROS_SV__
